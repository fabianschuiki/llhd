-- Copyright (c) 2014 Fabian Schuiki

-- §13.9  Reserved words
abs access after alias all and architecture array assert attribute begin block
body buffer bus case component configuration constant label disconnect downto
map else elsif end entity exit file for function generate generic group
guarded if impure in inertial inout is library linkage literal loop mod nand
new next nor not null of on open or others out package port postponed
procedural procedure process protected pure range record reference register
reject rem report return rol ror select severity shared signal sla sll sra srl
subtype then to transport type unaffected units until use variable wait when
while with xnor xor

ABS ACCESS AFTER ALIAS ALL AND ARCHITECTURE ARRAY ASSERT ATTRIBUTE BEGIN BLOCK
BODY BUFFER BUS CASE COMPONENT CONFIGURATION CONSTANT LABEL DISCONNECT DOWNTO
MAP ELSE ELSIF END ENTITY EXIT FILE FOR FUNCTION GENERATE GENERIC GROUP
GUARDED IF IMPURE IN INERTIAL INOUT IS LIBRARY LINKAGE LITERAL LOOP MOD NAND
NEW NEXT NOR NOT NULL OF ON OPEN OR OTHERS OUT PACKAGE PORT POSTPONED
PROCEDURAL PROCEDURE PROCESS PROTECTED PURE RANGE RECORD REFERENCE REGISTER
REJECT REM REPORT RETURN ROL ROR SELECT SEVERITY SHARED SIGNAL SLA SLL SRA SRL
SUBTYPE THEN TO TRANSPORT TYPE UNAFFECTED UNITS UNTIL USE VARIABLE WAIT WHEN
WHILE WITH XNOR XOR


-- Partial Reserved Words.
a b c d e f g i l m n o p r s t u v w x

ab ac af al an ar as at be bl bo bu ca co di do el en ex fi fo fu ge gr gu if im
in is la li lo ma mo na ne no nu of on op or ot ou pa po pr pu ra re ro se sh si
sl sr su th to tr ty un us va wa wh wi xn xo

acc aft ali arc arr ass att beg blo bod buf cas com con dis dow els ent exi fil
fun gen gro gua imp ine ino lab lib lin lit loo nan nex nul ope oth pac por pos
pro pur ran rec ref reg rej rep ret sel sev sha sig sub the tra typ una uni unt
var wai whe whi wit xno

acce afte alia arch arra asse attr begi bloc buff comp conf cons labe disc down
elsi enti func gene grou guar impu iner inou libr link lite othe pack post proc
prot rang reco refe regi reje repo retu sele seve shar sign subt tran unaf unit
unti vari whil

acces archi asser attri buffe compo confi const disco downt entit funct gener
gener guard impur inert libra linka liter other packa postp proce proce prote
recor refer regis rejec repor retur selec sever share signa subty trans unaff
varia

archit attrib compon config consta discon functi genera generi guarde inerti
librar linkag litera packag postpo proced proced proces protec refere regist
severi subtyp transp unaffe variab

archite attribu compone configu constan disconn functio generat inertia postpon
procedu procedu protect referen registe severit transpo unaffec variabl

architec attribut componen configur disconne postpone procedur procedur protecte
referenc transpor unaffect

architect configura disconnec procedura unaffecte

architectu configurat

architectur configurati
