library iee, whadup, iee.test, sup?;
