-- Copyright (c) 2014 Fabian Schuiki

a26_a42_t6_236_aSDf -- basic_identifier
\fsoue fja398' 0asdf?\ -- extended_identifier
